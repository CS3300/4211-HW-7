library verilog;
use verilog.vl_types.all;
entity hex_to_ASCII is
end hex_to_ASCII;
